<?xml version="1.0" encoding="utf-8"?>
<!-- Generator: Adobe Illustrator 16.0.0, SVG Export Plug-In . SVG Version: 6.00 Build 0)  -->
<!DOCTYPE svg PUBLIC "-//W3C//DTD SVG 1.1//EN" "http://www.w3.org/Graphics/SVG/1.1/DTD/svg11.dtd">
<svg version="1.1" id="Layer_1" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" x="0px" y="0px"
	 width="505.101px" height="165.036px" viewBox="0 0 505.101 165.036" enable-background="new 0 0 505.101 165.036"
	 xml:space="preserve">
<g>
	<path fill="#efddb8" d="M12.852,32.64c-0.137,1.09-1.906,3.742-5.304,7.956c-0.408,0.816-1.02,1.157-1.836,1.02
		c-1.09,0-2.11-0.408-3.06-1.224c-0.408-0.408-1.224-1.699-2.448-3.876C0.067,34.342,0,32.981,0,32.436
		c0.408-3.943,2.244-5.712,5.508-5.304c0.816,0.137,1.836,1.294,3.06,3.468c0.134,0.137,0.306,0.102,0.51-0.102
		c0.204-0.204,0.44-0.306,0.714-0.306c0.408,0,1.02,0.306,1.836,0.918C12.444,31.722,12.852,32.232,12.852,32.64z M150.552,26.112
		c-1.361,0.816-2.11,1.769-2.244,2.856c0,0.545,0.134,1.09,0.408,1.632c-0.682,0.274-1.565,0.886-2.652,1.836
		c0-0.134-0.07-0.338-0.204-0.612c-2.722,1.632-4.08,3.946-4.08,6.936c1.087-0.95,2.652-2.515,4.692-4.692l-0.204,1.02l1.224,0.204
		c0.408-0.134,0.679-0.204,0.816-0.204c-1.498,0-2.926,1.565-4.284,4.692c0,0.274,0.067,0.612,0.204,1.02
		c-2.856,4.896-4.284,7.889-4.284,8.976c0.408,0.137,0.816,0,1.224-0.408c0.408-1.087,2.244-3.535,5.508-7.344
		c-1.498,2.448-3.06,5.17-4.692,8.16c-3.13,6.12-4.762,9.929-4.896,11.424c0,0.274-0.239,0.851-0.714,1.734
		c-0.479,0.886-0.784,1.6-0.918,2.142c0,0.545,0.134,1.294,0.408,2.244l-0.612-0.408c0.271,0.274,0.408,0.612,0.408,1.02
		c0,0.274-0.204,0.612-0.612,1.02v0.408c-0.137,0.137-0.07,0.274,0.204,0.408l0.816-1.428c0.679,1.09,0.95,1.836,0.816,2.244
		c0,0.816-1.361,3.468-4.08,7.956c-0.137,0-0.204,0.408-0.204,1.224l-0.816-0.612v0.204c0,0.137,0.067,0.274,0.204,0.408
		c0.134,0.137,0.204,0.408,0.204,0.816c-0.137,0.408-1.02,2.652-2.652,6.732c-0.682-0.134-1.224-0.134-1.632,0
		c-0.137,0.545,0,0.816,0.408,0.816c0.271,0.137,0.612,0,1.02-0.408c-0.274,0.545-0.816,1.361-1.632,2.448
		c0.542,0.545,1.087,1.294,1.632,2.244l-11.628,26.112c-5.986,13.738-11.832,23.256-17.544,28.561c0,0.679-0.749,1.969-2.244,3.875
		c-0.682,0.271-1.632,0.883-2.856,1.836c-0.274,0-0.647-0.238-1.122-0.714c-0.478-0.478-0.851-0.714-1.122-0.714
		c-0.274,0-0.545,0.134-0.816,0.408c-0.274,0.271-0.545,0.408-0.816,0.408c-0.816,0-1.836-1.157-3.06-3.469
		c-0.682,0.271-1.02,0.746-1.02,1.429c0.134,0.679,0.134,1.224,0,1.632c-0.137-0.408-1.09-0.545-2.856-0.408
		c0.271,0.816,0.883,2.107,1.836,3.876c-6.936-2.993-10.2-4.488-9.792-4.488c-0.274,0-0.408,0.135-0.408,0.408
		c0,0.271-0.204,0.408-0.612,0.408c0.134,0,0.067-0.204-0.204-0.612c-3.946-1.224-6.802-1.836-8.568-1.836
		c-1.224-0.545-2.11-1.766-2.652-3.672c-0.137-0.271-0.545-0.541-1.224-0.816c-2.448-4.621-4.217-7.002-5.304-7.14
		c0-0.134,0.134-0.338,0.408-0.612l0.408-0.612c0.271-1.632-0.204-2.515-1.428-2.652c-0.953-0.134-2.04,1.09-3.264,3.672
		c0.134,0.274,0.204,0.682,0.204,1.224c-0.274,0-2.177,2.04-5.712,6.12c-3.538,4.08-5.849,6.051-6.936,5.917
		c0.408,0.134-0.478-0.408-2.652-1.633c-0.545,0-1.294-0.137-2.244-0.407c-0.953-0.274-1.702-0.408-2.244-0.408
		c-0.816,0.815-1.361,1.97-1.632,3.468c-0.408,0.679-1.361,0.883-2.856,0.612c-3.809-0.274-6.257-2.381-7.344-6.324l-3.672-4.08
		c-1.498-2.719-3.06-5.371-4.692-7.956c-1.769-3.535-2.926-6.391-3.468-8.568c-2.585-10.471-4.421-21.487-5.508-33.048l0.204-2.448
		c0-0.95-0.479-1.699-1.428-2.244c-0.408,8.705,0.338,16.661,2.244,23.868c-1.09-0.134-1.702-0.542-1.836-1.224
		c-0.545-1.766-1.02-3.943-1.428-6.528C0.95,95.609,0.746,86.362,1.836,76.296c0.271-2.99,1.291-5.642,3.06-7.956
		c-0.137,0.274-0.137-0.067,0-1.02c0.271,0.408,0.542,0.612,0.816,0.612l0.816-0.408c-0.408-0.271-0.816-0.95-1.224-2.04
		c0.542,0,0.95-0.134,1.224-0.408c0.271,0.816,0.679,1.906,1.224,3.264l0.816,0.204c0.271,0.274,0.475-0.271,0.612-1.632
		c-1.224-1.224-1.769-2.311-1.632-3.264c0.134,0,0.306-0.134,0.51-0.408c0.204-0.271,0.44-0.338,0.714-0.204
		c0.542,0,1.224,0.953,2.04,2.856c0.134-0.134,0.204-0.408,0.204-0.816c0.271-2.04-0.274-3.943-1.632-5.712
		c-0.137,0-0.306,0.035-0.51,0.102c-0.204,0.07-0.443,0.102-0.714,0.102c-0.408,0-1.02-0.848-1.836-2.55
		c-0.816-1.699-1.157-2.821-1.02-3.366c0-0.271,0.102-0.51,0.306-0.714s0.306-0.373,0.306-0.51H7.14
		c0.95,0.545,1.632,1.498,2.04,2.856c0.134,0.682,0,1.702-0.408,3.06c0.134,0.408,0.475,0.816,1.02,1.224
		c0.271-0.679,0.746-0.95,1.428-0.816c0.408,0.137,1.087,0.749,2.04,1.836c0.134-0.679,0.475-1.699,1.02-3.06
		c1.087,1.09,1.836,1.973,2.244,2.652c0.679,0.137,1.154,0.137,1.428,0c-2.722-4.759-4.013-7.819-3.876-9.18
		c0.134-0.95,0.883-2.244,2.244-3.876c1.358-1.632,2.515-2.378,3.468-2.244c0.679,0,1.562,0.612,2.652,1.836
		c1.087,1.224,1.562,2.177,1.428,2.856c0,0.545-0.306,1.428-0.918,2.652c-0.612,1.224-0.918,2.11-0.918,2.652
		c0.134,0.274,0.542,1.157,1.224,2.652c3.264-0.679,4.896-1.428,4.896-2.244c0,1.09-0.274-0.067-0.816-3.468
		c0.134,0,0.373-0.067,0.714-0.204c0.338-0.134,0.644-0.134,0.918,0c1.358,0.137,2.244,2.789,2.652,7.956
		c-0.545,13.056,0.542,27.406,3.264,43.044c0.271,0.408,0.679,1.157,1.224,2.244c0.271,0,0.475-0.134,0.612-0.408
		c0-0.134-0.137-0.338-0.408-0.612c1.224-1.495,1.699-2.515,1.428-3.06l0.816,1.02c0.542-0.679,0.883-1.224,1.02-1.632
		c-0.137-0.271-0.274-0.408-0.408-0.408c0.408-0.408,0.612-0.883,0.612-1.428c0.542-0.816,1.632-2.652,3.264-5.508
		c-0.137,0.274-0.545-0.067-1.224-1.02c0.542,0.137,0.883,0.274,1.02,0.408c0.271-0.271,0.679-0.746,1.224-1.428
		c0-0.134-0.07-0.338-0.204-0.612c0.816-1.087,1.358-2.311,1.632-3.672c1.358-1.495,2.174-2.786,2.448-3.876
		c0,0.137,0.134,0.274,0.408,0.408c0.816-0.542,1.358-1.495,1.632-2.856c0-0.542,0.067-1.428,0.204-2.652
		c0.816-0.271,1.326-1.052,1.53-2.346c0.204-1.291,0.985-2.346,2.346-3.162c1.358-0.816,2.244-1.428,2.652-1.836
		c0.134-4.351,1.02-8.906,2.652-13.668c0.408-1.224,1.428-2.582,3.06-4.08c1.632-1.495,2.99-2.174,4.08-2.04
		c1.224,0.137,2.378,1.294,3.468,3.468c0.408-0.271,1.087-0.338,2.04-0.204c-0.274-0.134,0.067-0.408,1.02-0.816l2.04-2.856
		l3.06,1.428c0.408,0,1.087-0.134,2.04-0.408c1.224,2.722,1.766,6.461,1.632,11.22L81.6,73.44c-0.137-0.408-0.274,0-0.408,1.224
		c0.134,0.274,0.271,0.408,0.408,0.408c0.408-0.408,0.679-0.95,0.816-1.632c0-0.408-0.137-1.087-0.408-2.04
		c0.271-0.271,0.679-0.338,1.224-0.204c0-0.679,0.134-1.632,0.408-2.856c0.271-1.224,0.475-2.174,0.612-2.856
		c0,0.545,0.204,1.294,0.612,2.244c0.134-0.408,0.612-1.632,1.428-3.672c0,0.137,0.067,0.204,0.204,0.204
		c0.271,0.137,0.542,0.137,0.816,0l-2.856,25.296c0-0.816-0.137-2.107-0.408-3.876c-0.408,0.545-0.682,1.361-0.816,2.448
		c-0.137,1.361,0,2.993,0.408,4.896c0.679-1.632,1.02-2.652,1.02-3.06l-0.612,16.932c-0.137,2.177-0.274,5.441-0.408,9.792
		c4.896-5.712,9.859-14.347,14.892-25.908c7.07-16.046,11.22-25.226,12.444-27.54c0.679-1.358,1.02-2.515,1.02-3.468
		c0.679-0.134,1.087-0.408,1.224-0.816c0-0.134-0.07-0.408-0.204-0.816c1.632-2.448,3.672-6.12,6.12-11.016
		c0,0.408,0.338,0.953,1.02,1.632c0.271,0,0.475,0,0.612,0c0.816-1.224,1.97-2.856,3.468-4.896c-0.953,3.264-2.652,6.732-5.1,10.404
		l0.408,1.02c-1.09,0.274-1.973,1.224-2.652,2.856c-0.274,0.682-0.408,1.294-0.408,1.836c-0.137,0.545,0,1.02,0.408,1.428
		c-0.137,0-0.408-0.271-0.816-0.816c-0.137,0.545-0.682,1.294-1.632,2.244v1.632c1.632-0.679,2.378-1.087,2.244-1.224
		c-0.545-0.408-0.816-0.746-0.816-1.02l0.816,0.204c-0.274,0,0.271-0.204,1.632-0.612c-0.408-0.542-0.478-0.816-0.204-0.816
		l0.204-0.204l0.204-0.816c0.134-0.271,1.699-2.856,4.692-7.752c0.408-0.95,0.338-1.495-0.204-1.632
		c0.408-0.134,0.883-0.612,1.428-1.428c0.408-1.495,1.291-3.672,2.652-6.528c1.632-1.495,3.194-3.264,4.692-5.304
		c0.408-0.408,1.766-2.107,4.08-5.1l2.04-2.448c-0.137,0.682-0.137,1.09,0,1.224c0.542-0.542,1.428-1.358,2.652-2.448l1.224-2.448
		c-0.137,0.137-0.07,0.341,0.204,0.612c0.408-0.542,0.816-1.154,1.224-1.836c0,1.632-0.545,3.197-1.632,4.692
		c0.134,0.137,0.338,0.204,0.612,0.204c0.408-0.408,1.495-1.495,3.264-3.264c-5.849,7.752-11.086,15.233-15.708,22.44
		c-0.408,0.816-0.545,1.632-0.408,2.448l13.056-17.544c0.542-0.816,1.154-1.699,1.836-2.652c-0.274,0-0.204,0.274,0.204,0.816
		c1.766-2.582,2.582-4.284,2.448-5.1c0.134,0,0.408,0.274,0.816,0.816c0.408-0.271,0.95-0.612,1.632-1.02
		c0.134-0.542,0.542-1.154,1.224-1.836V26.112z M29.376,18.768c-0.137,1.906-3.197,4.354-9.18,7.344
		c-1.498-1.358-2.856-2.107-4.08-2.244h-0.612c0,0.137-0.137,0.204-0.408,0.204c-3.809-0.408-5.374-3.806-4.692-10.2
		c0.408-3.535,1.766-5.167,4.08-4.896c0.816,0.137,1.428,0.341,1.836,0.612c2.99-4.351,5.234-6.458,6.732-6.324
		c1.903,0.274,3.331,1.498,4.284,3.672l1.836,5.916l-0.204,3.264c0,0.137,0.067,0.545,0.204,1.224
		C29.306,18.022,29.376,18.497,29.376,18.768z M17.544,39.984c-0.137,1.224-1.157,1.769-3.06,1.632
		c-1.09-0.134-2.04-1.087-2.856-2.856c0.679-0.816,1.495-1.154,2.448-1.02C16.524,37.877,17.678,38.626,17.544,39.984z M13.26,67.32
		h-0.612l-0.612,0.816l0.612,0.408L13.26,67.32z M13.464,85.272c0-1.766,0.067-4.147,0.204-7.14
		c-0.274-0.408-0.682-1.02-1.224-1.836l-0.204,1.836c0,0.953,0.271,1.973,0.816,3.06C12.374,82.961,12.511,84.322,13.464,85.272z
		 M13.668,62.628h-0.612l-0.408,1.02l0.612,0.204L13.668,62.628z M13.464,65.076V64.26h-0.408l-0.204,0.816H13.464z M18.36,80.784
		l-0.408-0.204l-0.408,0.816l0.408,0.408L18.36,80.784z M24.48,146.064l-1.02-0.204v-0.611l1.02,0.203V146.064z M27.744,74.052
		l0.204-2.856c-0.274-0.134-0.545-0.338-0.816-0.612c0,0.408-0.137,1.565-0.408,3.468l-0.408,0.204c0,0.274,0,0.612,0,1.02
		C26.45,75.005,26.928,74.597,27.744,74.052z M32.028,39.168c-2.993,1.361-4.217,2.04-3.672,2.04
		c-1.499-0.134-2.11-1.428-1.836-3.876c0.134-1.766,0.816-2.582,2.04-2.448c0.95,0.137,2.174,0.816,3.672,2.04L32.028,39.168z
		 M28.764,59.16v-0.816l-0.612-0.204v0.816L28.764,59.16z M51.408,22.032c-0.545,0.545-0.886,0.816-1.02,0.816
		c0.408,0-0.749-0.612-3.468-1.836c0-0.542,0.134-1.632,0.408-3.264c1.087,0.408,2.515,1.02,4.284,1.836L51.408,22.032z
		 M55.08,72.42l-0.408-0.204l-0.408,1.02l0.408,0.204L55.08,72.42z M66.096,56.712c0.271-2.174,0.271-3.398,0-3.672
		c-1.09,0.953-1.702,1.769-1.836,2.448c0,0.408,0.067,0.75,0.204,1.02v0.408c0.134,0,0.408-0.032,0.816-0.102
		C65.688,56.747,65.958,56.712,66.096,56.712z M78.744,121.584l1.632-26.52c0,0.408-0.102,1.122-0.306,2.142
		s-0.376,1.734-0.51,2.142L78.744,121.584z M80.988,93.228h-0.612l-0.408,1.02l0.612,0.204L80.988,93.228z M81.192,92.004H80.58
		l-0.408,1.02l0.408,0.204L81.192,92.004z M81.6,87.924c-0.274-1.358-0.341-2.311-0.204-2.856c-0.408,3.13-0.545,4.966-0.408,5.508
		C80.988,90.168,81.192,89.285,81.6,87.924z M82.008,82.212l0.408-4.08c-0.816,1.361-1.224,2.244-1.224,2.652
		C81.326,81.058,81.6,81.533,82.008,82.212z M82.824,76.704L82.212,76.5l-0.408,0.612l0.612,0.408L82.824,76.704z M83.028,111.18
		l0.408-3.06h-0.612l-0.408,3.06H83.028z M83.232,113.424l0.204-1.224h-0.612l-0.204,1.224H83.232z M83.436,117.096l-0.408,1.428
		l-0.408-0.204l0.408-1.224H83.436z M83.436,106.488l0.204-2.856h-0.612l-0.204,2.856H83.436z M83.64,100.164l0.204-1.224h-0.612
		l-0.204,1.224H83.64z M84.252,84.66l0.204-2.652h-0.612l-0.204,2.448L84.252,84.66z M103.836,91.188
		c-0.408,0-0.682-0.204-0.816-0.612c0.679-1.632,1.087-3.264,1.224-4.896c-0.816,1.361-1.836,3.264-3.06,5.712
		c0.271,0.816,0.338,1.428,0.204,1.836c0,0.545-0.341,1.09-1.02,1.632l-0.204,2.244c0.816-0.408,1.597-1.46,2.346-3.162
		C103.256,92.243,103.699,91.325,103.836,91.188z M103.02,147.493c-0.408,0.545-1.02,0.745-1.836,0.611
		c0.134,0.134,0.204,0.408,0.204,0.816C102.475,148.646,103.02,148.171,103.02,147.493z M104.448,146.268l-1.02,1.02l-0.204-0.408
		l0.816-1.02L104.448,146.268z M110.772,77.112c0-0.271-0.07-0.542-0.204-0.816c-0.137-0.271-0.204-0.475-0.204-0.612
		c-0.274,0-0.478,0.137-0.612,0.408c0.134,0.816-0.274,1.428-1.224,1.836c-0.408,1.906-1.361,4.15-2.856,6.732
		c0-1.087-0.07-1.903-0.204-2.448c0,0.408-0.172,0.918-0.51,1.53c-0.341,0.612-0.51,1.122-0.51,1.53l1.02-0.408
		c0.271,0.274,0.408,0.612,0.408,1.02C109.003,80.446,110.635,77.52,110.772,77.112z M106.692,81.192l0.204-1.02l-0.408,0.204
		c-0.274,0.137-0.408,0.274-0.408,0.408C106.08,81.058,106.284,81.192,106.692,81.192z M112.2,69.36l-0.408-0.204l-0.612,1.836
		h0.612L112.2,69.36z M114.24,70.176c0-0.134-0.035-0.373-0.102-0.714c-0.07-0.338-0.102-0.577-0.102-0.714
		c-0.274,0.408-0.682,0.953-1.224,1.632C113.22,70.109,113.695,70.042,114.24,70.176z M114.852,65.892h-0.612l-0.612,1.632
		l0.612,0.204L114.852,65.892z M126.684,57.12h-0.408l-0.408,1.02l0.204,0.408L126.684,57.12z M128.928,42.432l-0.204-0.612
		l-1.428,1.224l0.408,0.204L128.928,42.432z M128.316,89.556l-0.408-0.408l-0.408,0.204l0.408,0.612L128.316,89.556z M130.56,83.64
		c-0.682,0.953-1.157,1.632-1.428,2.04h0.612C130.152,84.73,130.423,84.048,130.56,83.64z M133.824,68.952l-0.612-0.204
		l-0.612,2.244h0.408L133.824,68.952z M134.028,21.42l-0.816,0.816l-0.408-0.204l0.612-1.02L134.028,21.42z M135.048,68.136v-1.428
		h-0.612v1.428H135.048z M137.7,73.644l-1.02,1.428l-0.408-0.204l1.02-1.224H137.7z M137.496,65.688l-1.02,0.204v-0.408l0.816-0.408
		L137.496,65.688z M140.556,18.564c-0.682,1.498-1.294,2.652-1.836,3.468c-0.137-0.271-0.204-0.612-0.204-1.02
		C138.516,20.604,139.195,19.788,140.556,18.564z M141.372,23.256h-0.612v-1.02h0.612V23.256z M143.412,16.116l-1.836,2.04
		l-0.408-0.408l1.836-2.04L143.412,16.116z M142.392,24.276l-1.224,1.02c0-0.542,0.338-1.291,1.02-2.244
		C142.188,23.597,142.255,24.005,142.392,24.276z"/>
	<path fill="#efddb8" d="M233.783,85.884c0,2.448-1.021,6.053-3.06,10.812c-0.816,2.314-1.973,5.986-3.468,11.016
		c-1.632,1.769-3.946,4.762-6.936,8.976l1.02-2.04c0.816-1.495,1.087-2.378,0.816-2.652c-1.09,1.498-2.585,3.946-4.488,7.344
		c-0.816,0.682-2.04,1.973-3.672,3.876c-0.816,1.499-1.973,3.672-3.468,6.528c-3.539,5.033-7.481,9.113-11.832,12.24
		c-7.481,5.578-12.444,8.364-14.892,8.364c-0.408,0-1.02-0.137-1.836-0.408c-0.816-0.274-1.361-0.408-1.632-0.408
		c-1.09,0-2.62,0.236-4.59,0.714c-1.973,0.476-3.503,0.715-4.59,0.715c-4.08,0-8.434-2.178-13.056-6.528l-4.08-0.816
		c-0.137,0.408-0.204,0.953-0.204,1.633c0,0.682,0.067,1.498,0.204,2.447c-1.361-1.766-3.197-4.08-5.508-6.936
		c-0.137-0.679-0.478-1.903-1.02-3.672c-0.408-0.271-0.816-0.542-1.224-0.816c-0.274-1.766-0.682-4.488-1.224-8.16
		c0.679-0.816,1.02-1.428,1.02-1.836c-1.361-3.127-2.244-5.779-2.652-7.956c0.408-0.408,0.408-4.08,0-11.016
		c1.224-9.926,3.739-19.718,7.548-29.376c1.495-4.214,4.418-8.635,8.772-13.26c4.622-5.438,8.772-8.568,12.444-9.384
		c0.542,0,3.127-1.087,7.752-3.264c-9.384,3.809-16.865,9.725-22.44,17.748c-0.137,0.137,0,0.408,0.408,0.816l1.02-0.816
		c-1.769,1.906-3.197,4.217-4.284,6.936l0.816,0.408c4.214-5.846,11.083-12.036,20.604-18.564c-0.408,0-1.565,0.341-3.468,1.02
		c8.702-5.167,15.434-7.682,20.196-7.548c-0.137,0-0.408,0.204-0.816,0.612c0.408,0.274,0.883,0.408,1.428,0.408
		c0.679,0,1.699-0.134,3.06-0.408c1.358-0.271,2.378-0.408,3.06-0.408c0.408,0,1.326,0.478,2.754,1.428
		c1.428,0.953,2.276,1.428,2.55,1.428c0.542,0,0.781-0.102,0.714-0.306c-0.07-0.204,0.032-0.306,0.306-0.306
		c0.408,0.137,0.985,0.581,1.734,1.326c0.746,0.749,2.754,2.958,6.018,6.63c0.542,1.224,1.903,2.856,4.08,4.896l0.816-0.816
		c-0.953-0.408-1.326-0.95-1.122-1.632c0.204-0.679,0.032-1.224-0.51-1.632c2.174,0,3.806,0.478,4.896,1.428
		c0.816-0.95,1.224-1.562,1.224-1.836c0.542,1.498,1.632,3.06,3.264,4.692c0.95,1.09,2.378,4.558,4.284,10.404
		c0,0.545,0.067,1.428,0.204,2.652c0.271,0.545,0.883,1.09,1.836,1.632C233.375,83.436,233.783,84.66,233.783,85.884z
		 M164.423,64.26l-2.652,2.856l-0.204-0.612l2.448-2.448L164.423,64.26z M167.687,62.22l-2.652,2.04l-0.204-0.816l2.448-1.836
		L167.687,62.22z M200.123,81.804c-1.361-2.04-2.177-3.602-2.448-4.692c-1.769,1.224-4.625,3.538-8.568,6.936
		c0.134-0.816,0.679-1.836,1.632-3.06c-6.257,7.752-10.812,16.39-13.668,25.908c-0.545-0.816-0.886-1.224-1.02-1.224
		c-0.953,0-1.871,1.632-2.754,4.896c-0.886,3.264-1.326,5.578-1.326,6.936c0,2.722,0.612,6.257,1.836,10.608
		c5.438-1.495,10.675-5.508,15.708-12.036c5.03-6.528,7.478-12.444,7.344-17.748c0.542,0.274,0.95-0.134,1.224-1.224l0.612-1.428
		c-1.09-0.408-2.244-0.883-3.468-1.428c0.134-0.679,0.204-1.224,0.204-1.632c0-1.358-2.177-2.582-6.528-3.672l5.1-0.204
		c0.679,0.274,1.632,0.886,2.856,1.836c0.134-0.408,0.338-0.883,0.612-1.428c-0.816,0-1.294-0.067-1.428-0.204
		c0.679-0.679,0.95-1.224,0.816-1.632c-0.545-0.408-1.294-0.95-2.244-1.632c2.04-0.679,3.398-1.562,4.08-2.652
		c-0.408-0.542-0.953-1.154-1.632-1.836c0.408,0,0.95,0.102,1.632,0.306C199.374,81.702,199.849,81.804,200.123,81.804z
		 M181.967,52.02h-1.224v-0.816h1.224V52.02z M190.739,52.224c-1.498,0.408-4.558,1.428-9.18,3.06h1.836
		C184.211,55.421,186.659,54.401,190.739,52.224z M184.619,51h-1.224v-0.816h1.224V51z M193.595,94.86h-1.02v-0.816h1.02V94.86z
		 M229.907,61.404h-0.816v-1.836h0.816V61.404z"/>
	<path fill="#efddb8" d="M230.109,38.76c1.903-0.816,3.398-1.428,4.488-1.836c0.134,1.632,0.204,2.722,0.204,3.264
		c-2.722,1.09-3.876,1.632-3.468,1.632c-0.137,0-0.478-0.204-1.02-0.612L230.109,38.76z M235.413,88.536l0.204-0.816l-0.204-2.04
		c1.495-3.535,2.856-5.371,4.08-5.508c0.95,0,1.836,0.612,2.652,1.836c0.271,0.816,0.678,1.565,1.223,2.244
		c0.271-0.134,0.68-0.204,1.225-0.204c1.357,0,2.107,1.02,2.244,3.06c0.135,3.946-0.953,5.916-3.264,5.916
		c-0.137,0-0.205-0.067-0.205-0.204l-0.406,0.204c-0.683,0-1.566,0.408-2.653,1.224c-3.538-2.582-5.304-4.147-5.304-4.692
		C235.006,89.285,235.14,88.944,235.413,88.536z M239.697,132.396l-2.244,7.548l0.408,0.204l2.448-7.752H239.697z M317.625,66.504
		c-0.406-1.632-0.406-2.582,0-2.856c-1.09-3.943-1.904-6.936-2.447-8.976c-1.906-1.495-3.131-2.311-3.672-2.448
		c-0.408,0.953-0.611,1.702-0.611,2.244h-0.408c-1.09-1.766-1.973-2.582-2.652-2.448l-2.447,1.428
		c-0.275-0.408-0.479-0.679-0.613-0.816c-2.721-1.632-4.488-2.378-5.303-2.244c-0.816,0-3.266,1.973-7.346,5.916
		c-0.682,0-1.223-0.271-1.631-0.816c0,0.682-0.137,1.157-0.408,1.428l-1.225,0.204c-0.273,0-0.375-0.102-0.305-0.306
		c0.066-0.204-0.035-0.306-0.307-0.306c-0.682,0-1.361,0.749-2.039,2.244v1.836c0,0.682-0.139,1.224-0.408,1.632
		c1.223-1.766,2.105-3.06,2.65-3.876l0.205,0.408c-5.033,8.842-9.113,15.574-12.24,20.196c-0.137-1.766-0.137-4.214,0-7.344
		c-0.137-0.134-0.203-0.271-0.203-0.408c0.406-3.672,0.406-6.732,0-9.18c-0.139,0-0.24,0.07-0.307,0.204
		c-0.07,0.137-0.24,0.204-0.51,0.204c-0.545,0-0.75-0.816-0.613-2.448l0.408-2.448c-2.992-3.264-5.236-4.488-6.73-3.672
		c2.719,1.361,4.01,2.448,3.875,3.264c1.088,0.274,1.699,1.157,1.836,2.652c0,0.545-0.07,0.953-0.203,1.224
		c-1.361-2.719-2.789-4.284-4.285-4.692c0,0.137,0.066,0.341,0.205,0.612c0.133,0.274,0.203,0.478,0.203,0.612l0.611-0.204
		c0.68,0,1.43,0.682,2.244,2.04l-1.631,0.816c-2.855-3.127-4.559-4.759-5.1-4.896c0.27-0.408,0.406-0.883,0.406-1.428
		c-2.313,1.498-4.486,2.448-6.527,2.856c-1.498,0.682-2.584,1.157-3.264,1.428c-0.137,0.545-0.203,1.02-0.203,1.428
		c-0.547,1.09-1.295,1.906-2.244,2.448c-1.225-0.408-2.178-0.679-2.857-0.816c0-0.134-0.203-0.067-0.611,0.204
		c0.271,0,0.408,0.137,0.408,0.408c-0.682,1.906-1.09,2.993-1.225,3.264c0.135-0.134,0.439-0.271,0.918-0.408
		c0.475-0.134,0.781-0.271,0.918-0.408c0.135,0.137,0.135,0.274,0,0.408c-1.498,1.906-2.244,3.06-2.244,3.468
		c-1.09,0.545-1.906,1.09-2.447,1.632l0.816-0.612c0.408,0.408,0.678,0.75,0.816,1.02c-0.139,0.274-0.139,0.612,0,1.02
		c0.541-1.495,0.949-2.377,1.223-2.652c0.271,0.545,0.205,1.02-0.203,1.428c0.678-0.134,0.949,0.478,0.816,1.836
		c0.949,4.217,1.494,6.598,1.631,7.14c0.135,0.816-0.137,2.722-0.816,5.712c0.135-0.134,0.408,0.137,0.816,0.816
		c-1.09,5.986-1.836,9.996-2.244,12.036c-1.77,9.521-3.061,15.504-3.875,17.952c-1.498,4.217-2.244,7.548-2.244,9.996
		c0,0.137-0.102,0.478-0.307,1.02c-0.203,0.545-0.307,0.953-0.307,1.224c0,0.545,0.135,0.816,0.408,0.816l5.713-17.748
		l-5.508,21.216c0.949-3.264,1.699-5.575,2.244-6.936c0,0.274-0.75,3.197-2.244,8.772c0-0.271,0.27-0.475,0.816-0.612l-2.449,6.12
		c-0.137-0.816,0.032-1.903,0.509-3.264c0.475-1.358,0.645-2.174,0.51-2.448c-0.953,3.401-1.498,5.374-1.631,5.916
		c0-0.134,0.067-0.271,0.204-0.408c0.134,0.816-0.682,4.15-2.448,9.996l-0.407-0.611c0.134,2.174-0.07,3.602-0.612,4.284
		c0.679-1.091,1.224-1.906,1.632-2.448c0.134,0.408,0.204,0.679,0.204,0.815c-0.137-1.09,0.271-2.518,1.224-4.284l0.408,0.613
		c0-0.135,0.067-0.338,0.204-0.613c0.134,0.816,0.032,1.767-0.306,2.856c-0.342,1.087-0.511,1.836-0.511,2.244
		c0.542-1.498,0.95-2.519,1.225-3.06c0.408,0.407,0.611,0.679,0.611,0.815c-0.682,1.766-1.02,3.061-1.02,3.876
		c1.631-3.264,2.514-5.033,2.653-5.304c8.293-21.895,12.443-32.911,12.443-33.048c2.582-8.293,4.758-16.045,6.527-23.256
		c0.951,0.953,1.428,1.294,1.428,1.02c-4.762,17.952-7.209,27.132-7.344,27.54c-3.264,12.24-6.801,22.032-10.607,29.376
		c0.408-0.274,0.611-0.204,0.611,0.204v1.224c0.543-1.769,1.291-3.264,2.244-4.488c0.271,0.138,0.338,0.275,0.205,0.408
		c-0.953,2.856-1.77,4.622-2.449,5.305c-1.906,3.806-3.129,6.799-3.672,8.976c0.816-1.632,1.428-2.789,1.836-3.468
		c0.135,0,0.135,0.134,0,0.408c0,0.134,0.135,0.204,0.408,0.204c0.271-0.138,1.496-2.586,3.672-7.345
		c3.398-7.344,5.168-11.149,5.305-11.424c0.133,0.137,0.203,0.408,0.203,0.816c0.135,0.954-1.428,4.966-4.691,12.037
		c0.816-1.091,1.563-2.04,2.244-2.856c0.133-0.408,0.271-0.545,0.408-0.408c0.408-0.273,0.746-0.273,1.02,0
		c-1.225,3.127-2.039,5.575-2.447,7.345c1.494-2.586,3.127-6.054,4.895-10.404l-0.611,0.612c0-0.408,0.408-1.496,1.225-3.265
		c0.271,0.274,0.408,0.479,0.408,0.612c0.27-2.174,0.611-3.739,1.02-4.692c0.408,0.408,0.475,0.749,0.203,1.02
		c3.127-5.983,4.693-10.471,4.693-13.464c1.357-2.174,2.039-3.806,2.039-4.896c0-0.408-0.203-0.746-0.611-1.02
		c0.541-0.408,0.883-0.679,1.02-0.816c0.135-1.224,0.408-1.97,0.816-2.244l-0.205-1.428c-0.273-0.542-0.203-1.154,0.205-1.836
		l0.611,0.408c0.543-1.495,0.951-2.582,1.225-3.264c-0.545,0.682-1.02,1.09-1.428,1.224c0-1.632,0.408-2.652,1.223-3.06
		c0.271,0.408,0.408,0.816,0.408,1.224c2.582-9.384,4.555-14.551,5.916-15.504l0.613,0.612c0.27-0.271,0.746-0.408,1.428-0.408
		c0.133-1.087,0.475-2.174,1.02-3.264c0.271,0.137,0.338,0.274,0.203,0.408c-0.273,1.632-0.682,3.06-1.223,4.284
		c-0.275-0.271-0.342-0.408-0.205-0.408c0.408,0.408,0.613,0.816,0.613,1.224c0,0.408-0.24,1.192-0.715,2.346
		c-0.479,1.157-0.58,2.008-0.307,2.55c1.359-2.719,2.174-4.214,2.449-4.488l0.408,0.408c-0.137,1.632-0.205,2.856-0.205,3.672
		c1.225-2.582,2.174-4.214,2.857-4.896l0.406,0.408c-0.273,0.816-0.34,1.769-0.203,2.856c0.949-1.224,1.633-2.244,2.039-3.06
		c0.68,0.953,1.359,1.428,2.041,1.428c0.541-0.95,0.883-1.699,1.02-2.244c0.271,0.274,0.338,1.157,0.205,2.652
		c2.039-3.943,3.264-6.254,3.672-6.936c0.133,0.137,0.27,0.478,0.408,1.02c1.766-3.127,2.785-4.963,3.059-5.508
		c0.135,0.274,0.205,1.02,0.205,2.244l0.611-0.612c0.271,0.274,0.543,0.408,0.816,0.408c0.271,0,1.563-1.903,3.875-5.712
		c2.313-3.806,3.604-5.712,3.877-5.712h0.816h0.408l0.408-1.632c0-1.087,0.338-1.632,1.02-1.632c0.408,0,1.223,0.239,2.447,0.714
		c1.225,0.478,2.041,0.714,2.449,0.714c0.27,0,0.611-0.271,1.02-0.816c-0.137-0.816-0.07-1.291,0.203-1.428
		c0.816,1.09,1.225,1.973,1.225,2.652c0.133-1.632,0.338-2.856,0.611-3.672c0.408,0.953,0.68,1.702,0.816,2.244l-0.611,0.816h1.631
		c-0.137-2.856-0.07-4.622,0.205-5.304c0.814-1.495,1.291-2.378,1.428-2.652C317.83,67.728,317.625,66.778,317.625,66.504z
		 M239.086,155.448l-0.408,1.225l0.408,0.204l0.407-1.429H239.086z M241.125,152.184l-0.407,1.02h0.407l0.408-0.815L241.125,152.184
		z M243.369,148.512l-0.406-0.204l2.242-7.548h0.408L243.369,148.512z M244.185,163.2l-0.816,1.632l0.613,0.204l0.611-1.632
		L244.185,163.2z M244.593,57.12c1.496-1.224,2.719-1.836,3.672-1.836c1.225-0.134,1.902,0.682,2.041,2.448
		c0.133,2.448-0.545,3.742-2.041,3.876c0.543,0-0.682-0.746-3.672-2.244V57.12z M246.021,161.772l-1.428,3.264h0.816l1.225-3.264
		H246.021z M245.818,139.944v-0.816h0.611v0.816H245.818z M246.837,125.052h-0.611l0.408-2.04h0.611L246.837,125.052z
		 M247.449,123.012h-0.408l0.816-5.1h0.613L247.449,123.012z M248.265,157.284l-0.816,0.816l0.408,0.408l0.816-0.816
		L248.265,157.284z M248.47,66.096h-0.613v1.02h0.613V66.096z M249.693,61.2c-0.545,0.545-1.02,1.361-1.428,2.448
		c0.271-0.95,0.746-1.562,1.428-1.836l0.816,0.408C250.101,61.678,249.828,61.337,249.693,61.2z M250.509,73.644l-0.816,1.224
		l0.613,0.408l0.611-1.428L250.509,73.644z M250.714,89.76h-0.613v1.02h0.613V89.76z M250.509,68.952v-1.02h0.611v1.02H250.509z
		 M251.529,85.884h-0.611l0.203,1.02h0.613L251.529,85.884z M252.345,66.3l-0.408-0.204l0.408-0.816l0.408,0.204L252.345,66.3z
		 M252.142,64.26c0.408-1.224,0.949-1.97,1.631-2.244l0.205,1.836C253.57,63.581,252.957,63.718,252.142,64.26z M252.55,68.34
		l-0.408-0.204l0.408-0.816h0.203L252.55,68.34z M252.957,117.708l-0.406-0.204l0.406-1.02l0.613,0.204L252.957,117.708z
		 M256.63,127.704l-0.408-0.204l0.408-2.04h0.611L256.63,127.704z M259.078,60.996c-0.137-1.358,1.02-2.107,3.469-2.244
		c0.949,0,1.766,0.478,2.447,1.428L259.078,60.996z M259.689,138.312v-0.816l0.613-0.204v0.816L259.689,138.312z M260.71,136.884
		l-0.408-0.204l1.02-3.06h0.408L260.71,136.884z M262.341,130.764v-0.816h0.611v0.816H262.341z M262.75,129.744l-0.203-0.816h0.611
		l0.203,0.816H262.75z M263.158,128.112v-1.224l0.611-0.204v1.224L263.158,128.112z M263.769,126.276l-0.203-1.224h0.611
		l0.205,1.224H263.769z M264.177,53.856c0-0.408,0.439-0.883,1.326-1.428c0.883-0.542,1.529-0.816,1.938-0.816
		c0.271,0,0.51,0.102,0.715,0.306c0.203,0.204,0.373,0.306,0.51,0.306c0.541-0.95,1.563-1.428,3.061-1.428
		c3.264-0.134,4.963,1.09,5.1,3.672c0.133,0.545,0,1.906-0.408,4.08L264.177,53.856z M264.789,89.964h-0.611l0.205-2.652h0.611
		L264.789,89.964z M264.382,124.032v-1.02h0.406v1.02H264.382z M265.402,90.168h-0.613l0.408-2.856h0.613L265.402,90.168z
		 M269.074,110.16l-0.408-0.204l0.203-0.816l0.613,0.204L269.074,110.16z M269.482,108.732h-0.408l0.408-1.836h0.611
		L269.482,108.732z M270.093,105.06l-0.408-0.204l0.613-1.428h0.611L270.093,105.06z M271.113,103.224l-0.408,0.204v-1.836
		l0.613-0.204L271.113,103.224z M271.521,74.256l-0.611-0.204l0.408-1.02h0.611L271.521,74.256z M271.521,77.52v-1.224h0.613v1.224
		H271.521z M272.337,75.48h-0.408v-2.244h0.611L272.337,75.48z M274.582,97.308l-0.408,1.836l0.408,0.204l0.611-1.836
		L274.582,97.308z M277.642,70.176h-0.613l0.205,0.816h0.611L277.642,70.176z M284.986,63.036l-0.408,1.02l0.408,0.204l0.408-1.224
		H284.986z M295.593,90.984l-1.225,1.02l0.408,0.408l1.225-1.224L295.593,90.984z M298.654,86.904l-0.408-0.204l0.408-0.816h0.408
		L298.654,86.904z M300.285,47.736c-0.406,0.545-0.885,0.816-1.428,0.816c1.766-0.134,2.652,0.341,2.652,1.428
		C301.509,48.756,301.101,48.01,300.285,47.736z M311.302,79.968c0-0.408-0.139-0.679-0.408-0.816c0,1.09-0.137,1.702-0.408,1.836
		h0.611C311.232,80.58,311.302,80.242,311.302,79.968z M312.525,69.564l-0.408-2.04h0.613l0.408,1.836L312.525,69.564z
		 M314.566,70.584c0.541,2.04,0.883,3.197,1.02,3.468c-1.225-2.04-1.906-3.194-2.039-3.468c0-0.271,0.066-0.612,0.203-1.02
		c0.135-0.408,0.203-0.679,0.203-0.816c0.543,0.408,0.951,0.612,1.225,0.612C315.177,69.497,314.974,69.905,314.566,70.584z
		 M318.033,75.276h-0.408V76.5h0.408V75.276z"/>
	<path fill="#efddb8" d="M455.324,100.368c-2.041-0.271-3.809,0.204-5.305,1.428c-0.273,0.545-0.748,1.157-1.428,1.836
		c-1.225,1.09-2.518,2.11-3.877,3.06c-1.631,1.498-2.381,2.856-2.242,4.08c-1.77,1.769-5.713,5.17-11.832,10.2
		c-0.139,0.137-0.07,0.341,0.203,0.612c1.902-0.816,3.33-1.699,4.283-2.652l1.43,1.428c0,0.545-0.07,0.749-0.205,0.612l0.816,0.204
		c1.494,0,3.602-1.224,6.324-3.672l-3.672,3.06c0.133,0.137,0.611,0.274,1.428,0.408c1.225,0,3.467-0.883,6.732-2.652l-0.205,1.428
		c-0.682,0.953-1.701,2.11-3.061,3.468c-1.498,0.408-3.264,1.632-5.303,3.672c0.541,0.274,1.428,0.137,2.652-0.408
		c-0.408,0.408-1.057,0.918-1.939,1.53c-0.885,0.612-1.529,1.122-1.938,1.53l1.02,1.224c-1.906-0.271-2.855,0.204-2.855,1.428v1.428
		c-0.273,0-1.225,0.408-2.855,1.224c0,0.408,0.475,0.612,1.428,0.612c-2.992,1.906-6.189,3.876-9.588,5.916l-1.225,1.225
		c0,0.273,0.135,0.816,0.408,1.632c0.135,0.545,0.066,1.091-0.203,1.632l-5.713,4.08c-2.447,1.903-4.42,2.856-5.916,2.856
		c-3.4-0.138-5.1,0.541-5.1,2.04l-5.508-0.204c-0.408,0.134-0.682,0.031-0.816-0.307c-0.137-0.341-0.342-0.58-0.611-0.714
		c-0.545,0-3.131,0.679-7.752,2.04c-2.857,0.816-5.916,1.154-9.18,1.021c-7.891-0.408-15.371-2.856-22.441-7.345
		c-0.137-0.273-0.408-0.682-0.816-1.224c-2.584-1.357-3.672-2.04-3.264-2.04c-0.545,0-0.885,0.07-1.02,0.204l0.408-0.408v-0.204
		h-0.611l-1.021-1.02c-0.682-0.816-1.361-1.154-2.039-1.021c0.271,0.545,0.816,1.428,1.631,2.652c-1.09-1.087-2.518-2.786-4.283-5.1
		c0-0.679-0.137-1.632-0.408-2.856c-1.09-2.311-2.518-5.983-4.283-11.016c-0.684,0.137-1.021,0.478-1.021,1.02
		c0,0.816,0.068,1.157,0.205,1.02c0-0.542-0.273-1.087-0.816-1.632l-0.611,0.612c-0.816,4.762-2.855,12.24-6.121,22.44
		c0.271,0.407-0.34,0.611-1.836,0.611c-0.273,0-0.748-0.273-1.428-0.815c-0.682-0.545-1.293-0.816-1.836-0.816
		c0-0.408,0.271-0.886,0.816-1.428c-0.137-0.271-0.887-0.746-2.244-1.429c-1.361,1.767-3.605,4.692-6.732,8.772l-1.428-1.632
		c0.949-1.224,1.428-1.973,1.428-2.244c0-0.545-0.479-1.428-1.428-2.652c-0.545,0.271-1.701,1.699-3.469,4.284
		c-0.814-1.224-1.768-2.722-2.855-4.487c-0.137,0.134-1.631,1.224-4.488,3.264c-1.223-2.448-1.836-4.146-1.836-5.1
		c0.135-0.95,0.613-1.766,1.428-2.448c-0.137-0.271-0.406-0.612-0.814-1.021h-1.021c-0.406,0-0.611,0.204-0.611,0.612v-1.429
		c0.816-0.541,1.633-1.494,2.447-2.855c1.225-3.535,2.244-9.247,3.061-17.136c0.271-0.408,0.543-1.224,0.816-2.448
		c0.135-0.271,0.203-1.562,0.203-3.876c0-2.174-0.137-3.739-0.406-4.692l1.836-1.428l5.303-46.716
		c2.311-20.263,4.623-35.7,6.936-46.308c0.543-2.174,2.174-7.07,4.896-14.688c0.271-3.127,0.338-0.883,0.205,6.732l-0.613,12.648
		c0.543,0,1.021-0.338,1.428-1.02c0.816-5.03,2.652-12.036,5.51-21.012c0.949,0.408,2.105,1.361,3.467,2.856
		c0.543-0.408,1.633-0.542,3.264-0.408c0.135,0,0.408,0.07,0.816,0.204c0.408,0.137,0.746,0.204,1.02,0.204
		c0.408,0,0.613-0.134,0.613-0.408c0-0.271,0.203-0.338,0.611-0.204c0.271,0,0.541,0.137,0.816,0.408
		c0.271,0.274,0.611,0.408,1.02,0.408c1.357,0.137,2.174-0.612,2.447-2.244l2.244,4.896c-0.137,3.401-0.07,5.304,0.205,5.712
		c0.133,1.361,0,3.672-0.408,6.936c0.271,0.953,0.541,2.11,0.816,3.468l-8.16,64.668c-0.275,2.585,0.816,5.17,3.264,7.752
		c0.271,0.682,1.291,2.314,3.061,4.896c9.518-7.615,19.176-20.059,28.967-37.332c0.543,0.545,1.496,1.294,2.857,2.244
		c-0.545,2.04-1.158,3.672-1.836,4.896l-0.205,1.428c0.816,0.137,1.633-0.338,2.447-1.428l1.633-2.652
		c0.271,0.274,0.541,0.408,0.816,0.408c-0.137,2.177-0.275,3.468-0.408,3.876c1.086-0.816,1.902-1.766,2.447-2.856l-7.547,15.096
		c-2.586,5.304-5.646,9.929-9.18,13.872c-0.408,0.408-1.734,1.804-3.979,4.182c-2.244,2.381-3.367,3.707-3.367,3.978
		c0-0.408,0.613,0.682,1.836,3.264c-0.545-0.542-1.293-1.358-2.242-2.448c-0.684,0.274-1.43,1.224-2.244,2.856l0.814,0.408
		c0.408,0.137-0.273,0.204-2.039,0.204c-0.682,0.274-0.887,0.545-0.611,0.816c-0.816,0.274-1.906,1.294-3.266,3.06
		c1.768,1.906,4.488,3.334,8.16,4.284c8.16,2.177,11.967,3.264,11.424,3.264c0.68,0,2.721,0,6.121,0l5.916-0.204l0.611,0.816
		c4.488,0.274,14.893-4.759,31.213-15.096c-2.178,1.632-6.461,4.488-12.852,8.568c0,0.953,0.475,1.428,1.428,1.428l14.482-7.956
		c9.385-5.304,15.027-7.886,16.934-7.752c0.27,0,0.408,0.07,0.408,0.204c0,0.137,0.203,0.204,0.611,0.204
		c0.541,0.137,1.664-0.102,3.365-0.714c1.699-0.612,2.889-0.918,3.57-0.918C452.126,99.281,453.283,99.689,455.324,100.368z
		 M333.943,10.608h-0.816l-1.02,5.712h0.613L333.943,10.608z M345.572,130.968h-0.816v-1.02h0.816V130.968z M347.611,131.172
		l-0.408-2.04l-0.814-0.204l0.406,2.04L347.611,131.172z M352.71,87.924l-2.039,1.632l-0.408-0.408l2.041-1.632L352.71,87.924z
		 M361.279,108.528l-0.408-0.408l-2.855,2.448l0.408,0.612L361.279,108.528z M359.035,11.016h-0.814v-1.02h0.814V11.016z
		 M359.648,91.8l-0.613-0.204l-0.408-1.428l0.613-0.204L359.648,91.8z M366.175,103.224l-0.408-0.204l-4.08,4.08l0.408,0.408
		L366.175,103.224z M363.931,145.86l-2.039-1.02l-0.205,0.611l2.041,1.021L363.931,145.86z M368.214,109.752h-1.223v-0.816h1.223
		V109.752z M372.091,63.24l-3.264,4.692l-0.613-0.408l3.266-4.896L372.091,63.24z M370.458,109.956l-0.203,0.612l-1.428-0.612
		v-0.612L370.458,109.956z M387.392,153.408c-4.896-0.682-8.027-1.157-9.385-1.428c-3.539-0.816-6.324-1.973-8.363-3.468h1.428
		c1.766,0.134,4.283,0.815,7.547,2.04c3.264,1.224,5.779,1.902,7.549,2.04C386.984,152.592,387.392,152.863,387.392,153.408z
		 M372.5,110.976l-0.205,0.612l-1.428-0.612v-0.612L372.5,110.976z M377.191,64.668l-1.225,1.632l-0.406-0.612l1.02-1.428
		L377.191,64.668z M378.21,61.2l-0.814,1.632l-0.613-0.204l0.816-1.428H378.21z M378.21,89.556l-0.406-0.408l-1.021,1.428
		l0.408,0.408L378.21,89.556z M395.755,68.748c-1.633,3.13-4.217,7.752-7.752,13.872c-2.314,2.856-5.645,7.14-9.996,12.852
		L395.755,68.748z M386.167,77.928h-0.611l-1.836,3.876l0.406,0.408L386.167,77.928z M439.207,108.936l-0.203-0.612l-2.652,1.224
		v0.612L439.207,108.936z M456.955,100.368l-1.223-0.204v-0.612l1.223,0.204V100.368z"/>
	<path fill="#efddb8" d="M472.666,48.96c-1.498,0.682-3.061,1.769-4.693,3.264c-0.137-0.271-0.408-0.408-0.814-0.408
		c-1.633,0-2.789,1.565-3.469,4.692c2.855-1.495,4.826-2.856,5.916-4.08c-0.682,0.545-1.02,1.09-1.02,1.632
		c0,0.408,0.27,0.816,0.814,1.224c-0.406,0.137-2.789,1.294-7.139,3.468l0.203,0.408l-1.02-0.204l-0.611,0.612
		c1.494,0.408,2.719,0.612,3.672,0.612c-0.275,0.137-0.887,0.612-1.836,1.428c-0.684-0.271-1.703,0.035-3.061,0.918
		c-1.361,0.886-1.973,1.667-1.836,2.346c-0.137,0.137-1.156,0.953-3.061,2.448c-0.137,0.274-0.07,0.408,0.205,0.408
		c-0.137,0-0.408,0.07-0.816,0.204c-0.408,0.137-0.682,0.204-0.816,0.204c0.135,0,0.408-0.134,0.816-0.408
		c-1.361-0.271-2.652,0-3.877,0.816l-1.836,1.224h-1.223c-0.139,0.137-0.205,0.274-0.205,0.408c0,0.274,0.135,0.545,0.408,0.816
		c-0.137-0.134-0.342-0.067-0.611,0.204c-0.275,0.274-0.545,0.408-0.816,0.408c-0.273,0-0.273-0.134,0-0.408
		c0.135-0.271,0-0.408-0.408-0.408c-0.816,0-2.855,0.816-6.119,2.448l-4.896,2.448l-3.264,1.02c-1.361,0.682-2.178,1.02-2.449,1.02
		l-0.814,0.612c-2.314,0.545-3.469,1.361-3.469,2.448c0,1.09,0.816,2.448,2.447,4.08c0.135,0.953,0.543,2.381,1.225,4.284
		c2.174,0.274,3.398,0.408,3.672,0.408c0.271,0,0.408-0.067,0.408-0.204c0-0.134,0.133-0.204,0.408-0.204
		c0.271,0,0.576,0.172,0.918,0.51c0.338,0.341,0.645,0.51,0.918,0.51c1.086,0,2.617,0.204,4.59,0.612
		c1.971,0.408,3.434,0.612,4.387,0.612c1.902,0.137,3.533,0.478,4.895,1.02l0.816-0.816c2.174,0.545,5.576,2.244,10.201,5.1
		l-0.408,0.204c0.27,0.816,1.02,1.906,2.244,3.264h1.02c0.408,0,0.541-0.067,0.408-0.204l2.447,2.652
		c-0.137,0.137-0.238,0.376-0.307,0.714c-0.068,0.341-0.172,0.58-0.305,0.714c4.488,2.993,6.732,4.829,6.732,5.508
		c0,0.545-0.104,1.396-0.307,2.55c-0.205,1.157-0.307,2.008-0.307,2.55c0,0.816,0.066,1.769,0.205,2.856
		c-0.408-0.271-0.75-0.408-1.021-0.408c0.271-0.679,0.408-1.428,0.408-2.244s-0.137-1.766-0.408-2.856
		c-0.953,5.578-1.768,9.658-2.447,12.24c-1.361,4.896-3.334,8.976-5.916,12.24c-0.137,0.274-0.479,0.816-1.02,1.632l0.408-0.612
		l-0.613-0.612c-0.408,0.545-1.02,1.224-1.836,2.04c0.135,0.137,0.338,0.274,0.613,0.408l1.02-0.612
		c-0.137,0.682-0.545,1.498-1.225,2.448c-1.09,0.545-2.652,1.499-4.691,2.856c-0.545-1.225-1.158-1.836-1.836-1.836
		c-0.137,0.137-1.158,0.479-3.061,1.02c-0.273,0.408-0.137,0.612,0.408,0.612c-0.682,1.361-1.564,2.04-2.652,2.04
		c-0.273,0-0.408-0.066-0.408-0.204c0-0.134-0.137-0.204-0.408-0.204c-0.273,0-0.646,0.172-1.121,0.51
		c-0.479,0.342-0.852,0.511-1.123,0.511c-0.137-0.271-0.406-0.612-0.814-1.021c-0.137,0.137-0.342,0.307-0.613,0.51
		c-0.273,0.205-0.477,0.377-0.611,0.511c0.68,0,1.154,0.137,1.428,0.407c-0.408,0-1.055-0.066-1.938-0.203
		c-0.887-0.135-1.529-0.204-1.938-0.204c0.408,0,0.746-0.134,1.02-0.408c-0.408-0.408-0.682-0.612-0.816-0.612
		c-0.545,0-1.02,0.204-1.428,0.612l1.02,1.224c-0.273-0.271-0.545-0.408-0.816-0.408l-0.408,0.613
		c0.408,0.407,0.746,0.611,1.021,0.611c-4.08,1.357-5.646,2.04-4.693,2.04l-1.223-0.408c-0.275,0-0.918,0.373-1.939,1.122
		c-1.02,0.746-1.666,1.122-1.938,1.122c-0.682,0-1.701,0.067-3.059,0.204c-1.361,0.134-2.383,0.204-3.061,0.204
		c-0.275,0-0.816-0.408-1.633-1.225c-0.137,0.271-0.07,0.612,0.205,1.021c-1.225,0.408-2.928,0.883-5.102,1.428
		c-9.791,1.225-16.727,1.836-20.807,1.836h-2.041c-0.816,0-2.447-0.478-4.895-1.428c-0.139,0-0.342-0.07-0.613-0.204h-1.02
		c-0.408,0-0.545,0.103-0.408,0.306c0.135,0.204,0.066,0.307-0.203,0.307c-0.275,0-0.613-0.138-1.021-0.408
		c-0.408-0.137-0.885-0.137-1.428,0c0.68,0.679,1.291,1.02,1.836,1.02h-0.816c-0.682,0.135-1.156,0.204-1.428,0.204
		c-0.273,0-0.646-0.238-1.121-0.714c-0.479-0.478-0.918-0.714-1.326-0.714c-0.682,0-1.02,0.338-1.02,1.021l-1.428-0.612
		c-0.953-0.408-1.43-0.749-1.43-1.021c0-0.137,0.068-0.273,0.205-0.407c-0.137-0.274-0.545-0.408-1.225-0.408h-0.816
		c-0.133,0.134-0.338,0.204-0.611,0.204c0.408,0-2.039-0.749-7.344-2.244c-1.633-0.545-8.568-1.77-20.809-3.672
		c0.408,0,0.613-0.271,0.613-0.816c3.809,1.361,6.664,2.04,8.566,2.04c0.684,0,1.158-0.134,1.43-0.407
		c-2.582-1.088-4.352-1.633-5.305-1.633c-0.271,0-0.439,0.07-0.51,0.204c-0.068,0.138-0.236,0.204-0.51,0.204
		c-0.135-0.271-0.613-0.612-1.428-1.02c-2.041-1.088-3.943-1.633-5.713-1.633c0-0.271,0.07-0.541,0.203-0.816
		c-1.357-1.086-3.193-2.718-5.508-4.896c-0.133-0.408,0-1.428,0.408-3.06c-0.271-0.134-0.611-0.612-1.02-1.428h1.225
		c-0.135,0,0,0.204,0.408,0.612l0.611-0.612c-0.408-0.134-1.563-0.816-3.469-2.04c-0.133-0.408-0.541-1.02-1.223-1.836
		c0.406-0.95,1.156-1.699,2.244-2.244c0-0.408-0.477-0.612-1.43-0.612c0.408-0.816,1.361-1.358,2.857-1.632
		c-0.135-1.358,0-2.174,0.408-2.448c1.631,0.408,4.217,0.886,7.752,1.428l0.611,0.612c0.408,0,1.09,0.274,2.039,0.816
		c0.275-0.271,0.408-0.679,0.408-1.224c2.314,1.224,4.014,1.836,5.102,1.836c0.682,0,1.02-0.475,1.02-1.428
		c0.137,0.274,0.408,0.408,0.816,0.408c0.545,0,0.814-0.271,0.814-0.816c0.684,0.408,1.566,0.886,2.652,1.428
		c4.08,0.816,7.006,1.224,8.771,1.224c0.275,0,0.479-0.134,0.613-0.408c0.137-0.271,0.34-0.408,0.611-0.408
		c0.273,0,0.51,0.239,0.715,0.714c0.203,0.478,0.443,0.714,0.713,0.714c0.816,0,2.008,0.172,3.57,0.51
		c1.563,0.341,2.754,0.51,3.57,0.51c5.438,0,11.15-0.204,17.137-0.612c-0.139-0.134-0.479-0.204-1.021-0.204
		c2.582-0.271,6.051-0.746,10.404-1.428c8.977-0.271,18.902-1.766,29.785-4.488c0.541-0.408,0.814-0.679,0.814-0.816
		c1.359-0.134,2.787-0.746,4.285-1.836c0-0.816-0.275-1.224-0.816-1.224h-0.816l1.225-0.612c-0.273-0.271-0.75-0.408-1.428-0.408
		c0.816-0.134,2.855-1.154,6.119-3.06l-7.955-1.836c1.631,0.545,2.922,0.816,3.875,0.816h5.1v-1.428
		c-4.486-0.542-9.588-1.495-15.299-2.856l-1.225,0.204c0.68,0.682,1.02,1.09,1.02,1.224c-1.359-0.542-2.518-0.816-3.467-0.816
		c0.133,0,0.338-0.134,0.611-0.408c-0.273-0.408-0.816-0.612-1.631-0.612c-0.684,0-1.225,0.137-1.633,0.408
		c-0.273,0.137-0.137,0.682,0.408,1.632c-0.682-0.134-2.789-1.428-6.324-3.876c-0.408,0.408-0.479,0.749-0.205,1.02
		c-0.682-0.408-1.359-0.612-2.039-0.612c-1.361,0-2.244,1.294-2.652,3.876c-0.816-0.408-1.631-0.612-2.447-0.612
		c-0.275,0-0.715,0.07-1.326,0.204c-0.611,0.137-1.055,0.204-1.326,0.204c-0.273,0.274-0.203,0.816,0.203,1.632
		c-1.631-0.134-2.926,0.137-3.875,0.816c0.271-0.816,0.066-1.766-0.611-2.856c-0.816,0.137-1.703,1.428-2.652,3.876
		c0.133-0.95,0.066-1.632-0.205-2.04h-1.02c-0.137,0.408-0.203,0.816-0.203,1.224c0,0.408,0.066,0.816,0.203,1.224
		c-0.545-0.134-1.156,0-1.836,0.408c-0.137-0.679-0.408-1.562-0.816-2.652c-0.545,0.682-1.428,1.294-2.652,1.836
		c0.271-0.542,0.816-1.087,1.633-1.632c0.135-1.087,0.408-2.244,0.816-3.468l-0.205-1.632c-0.273,0.274-0.408,0.545-0.408,0.816
		c0,0.137,0.068,0.274,0.205,0.408c-0.273,0.137-0.611,0.408-1.02,0.816c-0.684-0.542-0.953-1.224-0.816-2.04
		c0.133-1.087,0.133-1.97,0-2.652c-1.906,0.816-2.723,2.652-2.449,5.508c0-0.134-0.102-0.271-0.305-0.408
		c-0.205-0.134-0.307-0.338-0.307-0.612c0-0.816,0.949-2.856,2.855-6.12l-0.203-1.632c-0.408,0-0.816,0.545-1.225,1.632
		c-0.137-0.271-0.545-0.746-1.223-1.428c-0.953,0.408-1.43,1.09-1.43,2.04c-0.406-0.408-0.748-0.612-1.02-0.612h-0.611
		c-0.137,0.137-0.273,0.204-0.408,0.204c1.766-2.174,2.652-3.672,2.652-4.488c0-0.408-0.102-0.679-0.307-0.816
		c-0.203-0.134-0.307-0.338-0.307-0.612h-0.814c-1.09,0-1.975,0.682-2.652,2.04c-0.137,0-0.443-0.134-0.918-0.408
		c-0.479-0.271-0.852-0.408-1.123-0.408c0.408-3.806,4.215-12.444,11.424-25.908c2.721-2.856,5.916-7.003,9.59-12.444v1.428
		c1.494-1.495,3.672-3.468,6.527-5.916c2.174-1.357,3.602-2.311,4.283-2.856c1.904-1.495,2.924-2.719,3.061-3.672
		c2.039,0,5.846-1.562,11.424-4.692l7.957-4.488c3.941-1.357,6.186-2.719,6.73-4.08c0.135,0.137,0.408,0.204,0.816,0.204
		c0.68,0,2.174-0.746,4.488-2.244c-0.408-0.408-0.75-0.612-1.02-0.612l0.816-1.02c0.133,0,0.234,0.239,0.305,0.714
		c0.066,0.478,0.307,0.714,0.715,0.714s0.816-0.204,1.223-0.612c-0.273,0,0.068,0.478,1.021,1.428
		c0.678-0.271,1.699-0.746,3.059-1.428v2.448c-0.545-0.134-0.953-0.134-1.223,0v0.612L456.14,35.7
		c-0.408-0.134-0.682-0.204-0.814-0.204l-0.205,2.04c2.041,0,3.264-0.816,3.672-2.448c3.398-1.632,5.508-2.244,6.324-1.836
		c0,0.274-0.203,0.682-0.611,1.224c0.133,0.137,0.408,0.204,0.816,0.204c0.27-0.679,0.406-1.562,0.406-2.652l1.836,1.224
		c0.271,1.361,0.408,2.244,0.408,2.652c0,0.137-0.238,0.51-0.713,1.122c-0.479,0.612-0.715,1.122-0.715,1.53
		c0,0.274,0.205,0.886,0.613,1.836c0.133-0.271,0.203-0.746,0.203-1.428c0.135,0,0.338-0.134,0.611-0.408
		c0.271-0.271,0.613-0.408,1.021-0.408c0.27,0,0.338,0.137,0.203,0.408c-0.137,0.274-0.07,0.408,0.203,0.408
		c0.408,0,0.781-0.134,1.123-0.408c0.338-0.271,0.576-0.408,0.715-0.408c0,0.274-0.07,0.749-0.205,1.428V40.8
		c0.816,0.953,1.225,1.769,1.225,2.448c-0.137,0.408-0.682,2.448-1.633,6.12c0-0.816,0.135-1.291,0.408-1.428v-1.224
		c-0.137-0.271-0.342-0.408-0.611-0.408l-1.021,3.06c0.135,0.137,0.477,0.204,1.021,0.204c0.541,0,1.02-0.338,1.428-1.02
		C472.257,48.826,472.527,48.96,472.666,48.96z M338.025,134.844h-1.02v-0.612h1.02V134.844z M344.552,145.656l-1.836-0.407v-0.612
		l1.836,0.407V145.656z M358.425,146.676v-0.612h-1.225v0.612H358.425z M358.833,143.413v-0.613h-1.021v0.613H358.833z
		 M359.853,144.84v-0.612h-0.816v0.612H359.853z M361.281,145.249v-0.612h-1.225v0.612H361.281z M361.078,147.493v-0.613h-1.021
		v0.613H361.078z M361.281,144.228v-0.612h-0.816v0.612H361.281z M363.117,144.636v-0.612h-1.225v0.612H363.117z M364.953,146.064
		v-0.612l-2.447-0.408v0.612L364.953,146.064z M364.544,138.72v-0.612h-0.816v0.612H364.544z M365.361,144.84v-0.612h-1.633v0.612
		H365.361z M365.564,148.512V147.9l-1.836-0.407v0.611L365.564,148.512z M367.4,146.676v-0.612l-2.242-0.408v0.612L367.4,146.676z
		 M368.625,139.536v-0.612h-1.02v0.612H368.625z M369.644,146.676v-0.612h-1.428v0.612H369.644z M371.074,139.944v-0.612h-2.041
		v0.612H371.074z M371.48,147.084v-0.612h-1.02v0.612H371.48z M371.48,149.124v-0.611h-1.02v0.611H371.48z M372.91,149.124v-0.611
		h-1.021v0.611H372.91z M378.621,146.676v-0.612l-5.916-0.408v0.612L378.621,146.676z M378.212,147.696v-0.611l-5.508-0.205v0.613
		L378.212,147.696z M374.949,149.532v-0.611h-2.039v0.611H374.949z M379.64,150.348v-0.612l-3.875-0.815v0.611L379.64,150.348z
		 M380.662,149.94v-0.612h-0.816v0.612H380.662z M381.884,153l-1.631-0.816l-0.205,0.612l1.633,0.815L381.884,153z M383.72,147.084
		v-0.612h-1.836v0.612H383.72z M386.169,143.004v-0.612h-3.061v0.612H386.169z M386.169,150.348v-0.612h-2.449v0.612H386.169z
		 M425.132,150.96c-0.545,0-1.396-0.07-2.549-0.204c-1.158-0.138-2.008-0.204-2.551-0.204c-0.273,0-0.545,0.169-0.816,0.51
		c-0.273,0.338-0.545,0.51-0.816,0.51c-0.273,0-0.545-0.102-0.814-0.306c-0.275-0.204-0.479-0.306-0.613-0.306
		c-1.631,0-3.197,0.338-4.691,1.02l-0.816-0.816c-1.09,0.135-2.721,0.542-4.895,1.225c0.27-0.274,0.406-0.545,0.406-0.816h-2.447
		c0,0.271-0.07,0.542-0.203,0.816c-0.408-0.408-0.816-0.612-1.225-0.612c0.408,0.408,0.541,0.679,0.408,0.816
		c-1.09-0.274-2.041-0.408-2.855-0.408c0.678,0,0.814,0.134,0.406,0.408h-1.02c-0.408-0.408-1.225-0.612-2.447-0.612h-5.1
		c-0.408,0.134-1.836,0.204-4.285,0.204h-2.855c0.541,0,1.393,0.306,2.551,0.918c1.152,0.612,1.867,0.918,2.141,0.918
		c0.271,0,0.68-0.102,1.225-0.306c0.541-0.204,0.949-0.307,1.225-0.307c0.27,0,0.27,0.134,0,0.408
		c-0.139,0.134-0.07,0.204,0.203,0.204c0.541,0,1.291-0.102,2.244-0.306c0.949-0.204,1.633-0.307,2.039-0.307
		c0.543,0.408,0.885,0.612,1.021,0.612c3.396,0,5.779-0.137,7.139-0.408c0-0.682,0.068-1.09,0.205-1.224
		c0.133,0,0.203,0.169,0.203,0.51c0,0.338,0.205,0.51,0.613,0.51c0.541,0,0.744-0.137,0.611-0.407l0.611,0.815
		c2.857,0,5.576-0.408,8.16-1.224c-0.273,0.271-0.07,0.408,0.613,0.408c1.223,0,2.58-0.408,4.08-1.225
		c0,0.271,0.475-0.07,1.428-1.02l0.203,0.611c0.135,0.408,0.408,0.612,0.816,0.612c0.271,0,0.713-0.172,1.326-0.51
		C424.623,151.129,424.996,150.96,425.132,150.96z M387.597,147.084v-0.612h-2.041v0.612H387.597z M388.414,150.144l-1.43-0.408
		v0.408l1.225,0.408L388.414,150.144z M390.861,126.888h-1.02v-0.612h1.02V126.888z M391.064,80.172l-0.611,1.428l-0.408-0.204
		l0.408-1.224H391.064z M392.085,77.316l-0.816,2.448l-0.611-0.204l0.814-2.244H392.085z M392.085,98.124v-1.02h-0.613v1.02H392.085
		z M394.125,150.348v-0.612h-2.039v0.612H394.125z M394.125,99.96l-0.203-0.612l-0.816,0.408v0.612L394.125,99.96z M400.041,147.493
		v-0.613h-5.1v0.613H400.041z M396.166,150.348v-0.612h-1.021v0.612H396.166z M397.593,150.348v-0.612h-1.02v0.612H397.593z
		 M399.429,128.316v-0.612h-2.449v0.612H399.429z M399.429,150.348v-0.612h-1.02v0.612H399.429z M403.304,128.316v-0.612
		l-3.467-0.204v0.612L403.304,128.316z M401.876,150.348v-0.612h-2.039v0.612H401.876z M400.857,151.368v-0.611h-1.02v0.611H400.857
		z M401.673,157.284l-0.205,0.612l-1.02-0.612l0.205-0.407L401.673,157.284z M404.121,156.468h-2.039v-0.816h2.039V156.468z
		 M403.304,150.348v-0.612h-0.814v0.612H403.304z M404.937,59.568l-1.225,1.224l-0.408-0.408l1.225-1.224L404.937,59.568z
		 M405.957,151.368v-0.611h-2.447v0.611H405.957z M405.548,150.348v-0.612h-1.631v0.612H405.548z M409.017,147.084v-0.612h-1.225
		v0.612H409.017z M410.242,156.468c-0.816,0-1.361,0.134-1.633,0.408l0.816-1.021C409.558,155.99,409.833,156.194,410.242,156.468z
		 M409.628,145.86l-0.611-0.408l-0.205,0.408l0.408,0.408L409.628,145.86z M418.4,155.04c-1.904,0.408-3.672,0.612-5.303,0.612
		c2.582-0.815,3.672-1.224,3.264-1.224C417.041,154.428,417.718,154.632,418.4,155.04z M415.953,150.552v-0.612h-1.428v0.612
		H415.953z M416.361,149.532v-0.611h-1.428v0.611H416.361z M417.38,145.656v-0.612h-1.428v0.612H417.38z M422.48,154.224h-1.836
		v-0.612h1.836V154.224z M423.91,153.612h-1.43V153h1.43V153.612z M426.765,150.348h-2.652c0.949,0,1.699,0.271,2.244,0.815
		C426.357,151.027,426.492,150.756,426.765,150.348z M430.232,151.368v-0.611h-0.814v0.611H430.232z M432.476,148.92v-0.612h-1.02
		v0.612H432.476z M433.089,147.696v-0.611h-1.225v0.611H433.089z M433.292,149.532l-0.203-0.611l-1.225,0.407v0.612L433.292,149.532
		z M434.517,147.493v-0.613h-1.225v0.613H434.517z M435.333,111.588h-1.021v-0.612h1.021V111.588z M438.597,117.096l-1.02,0.408
		v-0.408l0.814-0.408L438.597,117.096z M440.025,149.736l-1.225,0.816l-0.203-0.408l1.225-0.816L440.025,149.736z M442.064,146.064
		v-0.612h-1.223v0.612H442.064z M444.921,147.493h-0.816v-0.613h0.816V147.493z M448.593,138.108v-0.612h-1.02v0.612H448.593z
		 M448.593,144.024l-0.205-0.408l-0.814,0.408v0.408L448.593,144.024z M451.246,136.884l-0.205-0.408l-2.244,0.612v0.612
		L451.246,136.884z M450.224,150.144l-1.223,0.408v-0.408l1.02-0.408L450.224,150.144z M457.57,96.696
		c-0.547-1.087-3.197-2.311-7.957-3.672c-0.137,0.137-0.203,0.749-0.203,1.836C452.398,95.134,455.121,95.746,457.57,96.696z
		 M450.429,139.128v-0.612h-1.02v0.612H450.429z M458.384,139.536c-1.631,0.137-2.926,1.157-3.875,3.06
		c-0.137-0.271-0.408-0.408-0.816-0.408c0,0.273,0.135,0.682,0.408,1.225C456.14,142.461,457.57,141.168,458.384,139.536z
		 M460.22,65.484l-4.283,1.836v-0.408l4.08-2.04L460.22,65.484z M458.384,97.716l-2.039-0.816v0.612l1.836,0.612L458.384,97.716z
		 M459.201,100.572l-1.225-1.836l-0.406,0.408l1.223,1.632L459.201,100.572z M458.589,147.084h-0.816v-0.612h0.816V147.084z
		 M461.853,100.572c-1.225,0.682-1.77,1.224-1.633,1.632c0.543,0.545,0.951,0.816,1.225,0.816c0-0.271,0.066-0.679,0.203-1.224
		C461.783,101.254,461.853,100.846,461.853,100.572z M461.242,65.28h-1.021v-0.612h1.021V65.28z M462.669,137.496l-1.633,1.632
		l-0.203-0.408l1.631-1.632L462.669,137.496z M462.669,42.432l-0.205-0.408l-1.223,0.816l0.203,0.408L462.669,42.432z
		 M462.669,62.628l-1.021,0.816l-0.406-0.612l1.223-0.816L462.669,62.628z M464.097,56.916h-1.428l-0.613,0.816
		C462.873,57.732,463.552,57.461,464.097,56.916z M464.505,103.02c-0.545-0.408-1.225-1.087-2.041-2.04
		c0.135,0.274,0.205,0.545,0.205,0.816c0,0.408-0.137,0.749-0.408,1.02c1.086,1.09,1.631,1.565,1.631,1.428
		C463.892,103.702,464.097,103.294,464.505,103.02z M466.544,39.372c-0.682-0.134-1.428-0.542-2.244-1.224
		c-0.273-0.271-0.479-0.408-0.611-0.408v1.224c-0.137,0.545-0.205,0.886-0.205,1.02c0.135-0.134,0.271-0.338,0.408-0.612
		c0.135-0.271,0.271-0.475,0.408-0.612c0.271,0.816,0.135,1.565-0.408,2.244l-0.814,1.02
		C464.98,41.753,466.136,40.87,466.544,39.372z M464.708,59.364h-1.225v-0.612h1.225V59.364z M466.341,58.548l-1.02,0.612v-0.612
		l0.814-0.408L466.341,58.548z M466.75,134.64h-0.613l-0.408-0.816l0.613-0.204L466.75,134.64z M467.769,42.432l-0.408-0.408
		l-0.816,0.816l0.408,0.408L467.769,42.432z M468.177,49.572v-1.224h-0.613v1.224H468.177z M470.216,44.064v-4.08
		c-0.273-0.271-0.748-0.408-1.428-0.408c0,0.274-0.137,0.612-0.408,1.02c-0.273,0.408-0.408,0.816-0.408,1.224l0.613,0.612v2.856
		C468.994,45.017,469.535,44.609,470.216,44.064z M469.605,46.104l-0.205-0.612l-1.223,0.408v0.612L469.605,46.104z
		 M470.013,118.524H469.4v-1.02h0.613V118.524z M472.257,22.236l-0.816,0.816h-1.836v-2.448l1.428-1.428
		C471.304,19.313,471.712,20.333,472.257,22.236z M471.033,119.544h-0.611l-0.408-0.816l0.611-0.204L471.033,119.544z
		 M487.761,33.456c0,0.953-0.682,2.177-2.041,3.672l-2.447,2.04c-0.273-0.271-0.887-1.087-1.836-2.448
		c-0.408,0.274-1.428,0.07-3.061-0.612c0.816-0.542,1.291-1.087,1.428-1.632c-2.447-0.679-4.15-2.786-5.1-6.324l-1.428,1.428
		l-2.447-2.448c1.086-1.766,1.902-2.652,2.447-2.652l0.611,0.816c0.135-0.816,0.477-1.903,1.021-3.264
		c1.631-2.448,3.672-3.672,6.119-3.672c0.271,0,0.949,0.204,2.041,0.612c1.086,0.408,1.902,0.612,2.447,0.612
		c0.133,0.545,0.066,1.157-0.205,1.836c1.633,1.632,2.449,2.926,2.449,3.876c0,0.545-0.816,2.244-2.449,5.1
		C486.945,31.349,487.761,32.369,487.761,33.456z M473.48,124.44l-0.406,1.428l-0.408-0.204l0.408-1.224H473.48z M503.673,43.248
		c-1.906,1.361-4.83,3.264-8.773,5.712c-1.09,0.953-2.584,2.244-4.486,3.876c-0.139,0-0.408-0.134-0.816-0.408
		C491.636,49.301,496.33,46.241,503.673,43.248z M505.101,37.944c0,0.274-0.07,0.612-0.205,1.02
		c-0.137,0.408-0.203,0.749-0.203,1.02c-0.682-0.134-1.361,0-2.039,0.408c-0.547-0.679-0.816-1.087-0.816-1.224
		c0-0.271,0.133-0.781,0.408-1.53c0.27-0.746,0.408-1.256,0.408-1.53c0.541-0.134,1.357-0.134,2.447,0V37.944z"/>
</g>
</svg>
